module top_module (
	input clk,
	input L,
	input r_in,
	input q_in,
	output reg Q);

DFFMUX mod_inst1

endmodule

module DFFMUX (
	input clk,
	input L,
	input r_in,
	input q_in,
	output reg Q);
	
always @(posedge clk) begin
if (r_in) 
end
	
endmodule